module example(a,b,c);

input a;
input b;
output c;
assign c = a == b; 
initial begin
$display("hello ");

end
endmodule
