module adder(input [0:7] a,
	     input [0:7] b,
	     output [0:7] c);

assign c = a + b;
endmodule
